----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:33:23 04/14/2019 
-- Design Name: 
-- Module Name:    mux2x1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux2x1 is
  port(
    sw : in std_logic;
    x : in std_logic_vector(1 downto 0);
    y : out std_logic
  );
end mux2x1;

architecture behavior of mux2x1 is
  begin
    process(sw, x)
    begin
        if(sw = '0') then
          y <= x(0);
        elsif(sw = '1') then
          y <= x(1);
        else
          y <= 'Z';
        end if;
    end process;
end behavior;

